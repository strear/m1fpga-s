module indicator(
    input clk,
    input [1:0] mode,
    output [7:0] disp_an,
    output [6:0] disp_o
);

    reg [23:0] interval_c = 0;
    reg [7:0] t = 0;

    reg [6:0] disp [0:7];

    reg [2:0] sel = 0;
    assign disp_o = disp[sel];
    assign disp_an = sel == 7 ? 8'b01111111 : sel == 6 ? 8'b10111111
                   : sel == 5 ? 8'b11011111 : sel == 4 ? 8'b11101111
                   : sel == 3 ? 8'b11110111 : sel == 2 ? 8'b11111011
                   : sel == 1 ? 8'b11111101 : 8'b11111110;

    wire [7:0] f, g;
    assign f = ((t % 16 - 8) * (t % 16 - 8) * (t % 16 - 8) + 562) / 125;
    assign g = (((t + 8) % 16 - 8) * ((t + 8) % 16 - 8) * ((t + 8) % 16 - 8) + 562) / 125;

    always @(posedge clk) begin
        
        if (interval_c % 131072 == 0) sel = sel + 1;

        if (interval_c == 0) t = t + 1;

        case(mode)
            0: begin
                {disp[7], disp[6], disp[5], disp[4], disp[3], disp[2], disp[1], disp[0]} <= {
                    f == 0 ? 7'b0100011 : g == 0 ? 7'b0011100 : 7'b1111111,
                    f == 1 ? 7'b0011100 : g == 1 ? 7'b0100011 : 7'b1111111,
                    f == 2 ? 7'b0011100 : g == 2 ? 7'b0100011 : 7'b1111111,
                    f == 3 ? 7'b0011100 : g == 3 ? 7'b0100011 : 7'b1111111,
                    f == 4 ? 7'b0011100 : g == 4 ? 7'b0100011 : 7'b1111111,
                    f == 5 ? 7'b0011100 : g == 5 ? 7'b0100011 : 7'b1111111,
                    f == 6 ? 7'b0011100 : g == 6 ? 7'b0100011 : 7'b1111111,
                    f == 7 ? 7'b0100011 : g == 7 ? 7'b0011100 : 7'b1111111
                };
            end

            1: begin
                {disp[7], disp[6], disp[5], disp[4], disp[3], disp[2], disp[1], disp[0]} <= {
                      (t + 0) % 6 == 0 || (t + 0) % 6 == 1 ? 7'b1110111
                    : (t + 0) % 6 == 3 || (t + 0) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 1) % 6 == 0 || (t + 1) % 6 == 1 ? 7'b1110111
                    : (t + 1) % 6 == 3 || (t + 1) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 2) % 6 == 0 || (t + 2) % 6 == 1 ? 7'b1110111
                    : (t + 2) % 6 == 3 || (t + 2) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 3) % 6 == 0 || (t + 3) % 6 == 1 ? 7'b1110111
                    : (t + 3) % 6 == 3 || (t + 3) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 4) % 6 == 0 || (t + 4) % 6 == 1 ? 7'b1110111
                    : (t + 4) % 6 == 3 || (t + 4) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 5) % 6 == 0 || (t + 5) % 6 == 1 ? 7'b1110111
                    : (t + 5) % 6 == 3 || (t + 5) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 6) % 6 == 0 || (t + 6) % 6 == 1 ? 7'b1110111
                    : (t + 6) % 6 == 3 || (t + 6) % 6 == 4 ? 7'b1111110 : 7'b0111111,
                      (t + 7) % 6 == 0 || (t + 7) % 6 == 1 ? 7'b1110111
                    : (t + 7) % 6 == 3 || (t + 7) % 6 == 4 ? 7'b1111110 : 7'b0111111
                };
            end

            2: begin
                {disp[7], disp[6], disp[5], disp[4], disp[3], disp[2], disp[1], disp[0]} <= {
                    7'b1111111, 7'b1111111, 7'b1111001, 7'b1000000,
                    7'b0000110, 7'b0101111, 7'b0101111, 7'b1111111
                };
            end
        endcase
        
        interval_c = interval_c + 1;
    end
    
endmodule